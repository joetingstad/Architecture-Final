------------------------------------------------------------------------------------
---- Company: 
---- Engineer: 
---- 
---- Create Date: 04/21/2020 03:52:36 PM
---- Design Name: 
---- Module Name: generic_shifter - Behavioral
---- Project Name: 
---- Target Devices: 
---- Tool Versions: 
---- Description: 
---- 
---- Dependencies: 
---- 
---- Revision:
---- Revision 0.01 - File Created
---- Additional Comments:
---- 
------------------------------------------------------------------------------------


--library IEEE;
--use IEEE.STD_LOGIC_1164.ALL;

---- Uncomment the following library declaration if using
---- arithmetic functions with Signed or Unsigned values
----use IEEE.NUMERIC_STD.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx leaf cells in this code.
----library UNISIM;
----use UNISIM.VComponents.all;

--entity generic_shifter is
--    generic(width: integer := 32);
--    Port (shamt: in STD_LOGIC_VECTOR(9 downto 0);
--          a: in STD_LOGIC_VECTOR(width-1 downto 0);
--          output: out STD_LOGIC_VECTOR(width-1 downto 0));
--end generic_shifter;

--architecture Behavioral of generic_shifter is
----signal shamt
--begin
--    output <= 

--end Behavioral;
